* C:\Users\AWAIS SADDIQUI\Desktop\my cpp\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Tue Apr 12 11:44:19 2022



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
