* C:\Users\AWAIS SADDIQUI\Desktop\Playground\C&S -1\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Tue Apr 12 12:08:30 2022



** Analysis setup **
.DC LIN V_V1 1 50 1 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
